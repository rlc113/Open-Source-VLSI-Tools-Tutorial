module counter (clk,
    rst,
    out);
 input clk;
 input rst;
 output [28:0] out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_1 _077_ (.A(net2),
    .Y(_000_));
 sky130_fd_sc_hd__xor2_1 _078_ (.A(_057_),
    .B(net23),
    .X(_012_));
 sky130_fd_sc_hd__nand2_1 _079_ (.A(net23),
    .B(_056_),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _080_ (.A(net24),
    .B(_032_),
    .Y(_013_));
 sky130_fd_sc_hd__nand3_1 _081_ (.A(_057_),
    .B(net23),
    .C(net24),
    .Y(_033_));
 sky130_fd_sc_hd__xnor2_1 _082_ (.A(net25),
    .B(_033_),
    .Y(_014_));
 sky130_fd_sc_hd__nand4_1 _083_ (.A(net23),
    .B(net24),
    .C(net25),
    .D(_056_),
    .Y(_034_));
 sky130_fd_sc_hd__xnor2_1 _084_ (.A(net26),
    .B(_034_),
    .Y(_015_));
 sky130_fd_sc_hd__xor2_1 _085_ (.A(_060_),
    .B(net28),
    .X(_016_));
 sky130_fd_sc_hd__inv_1 _086_ (.A(net29),
    .Y(_035_));
 sky130_fd_sc_hd__nand4_2 _087_ (.A(net25),
    .B(net26),
    .C(net28),
    .D(net27),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _088_ (.A(_033_),
    .B(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__xnor2_1 _089_ (.A(_035_),
    .B(_037_),
    .Y(_017_));
 sky130_fd_sc_hd__nand3_1 _090_ (.A(net23),
    .B(net24),
    .C(_056_),
    .Y(_038_));
 sky130_fd_sc_hd__nor3_2 _091_ (.A(_035_),
    .B(_038_),
    .C(_036_),
    .Y(_039_));
 sky130_fd_sc_hd__xor2_1 _092_ (.A(net30),
    .B(_039_),
    .X(_018_));
 sky130_fd_sc_hd__xor2_1 _093_ (.A(_062_),
    .B(net4),
    .X(_001_));
 sky130_fd_sc_hd__xor2_1 _094_ (.A(_064_),
    .B(net6),
    .X(_002_));
 sky130_fd_sc_hd__xor2_1 _095_ (.A(_066_),
    .B(net8),
    .X(_003_));
 sky130_fd_sc_hd__nand4_1 _096_ (.A(net6),
    .B(net5),
    .C(net8),
    .D(net7),
    .Y(_040_));
 sky130_fd_sc_hd__nand3_1 _097_ (.A(net30),
    .B(net4),
    .C(net3),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_1 _098_ (.A(_040_),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__nor3_1 _099_ (.A(_035_),
    .B(_033_),
    .C(_036_),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _100_ (.A(_042_),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__xnor2_1 _101_ (.A(net9),
    .B(_044_),
    .Y(_004_));
 sky130_fd_sc_hd__nand3_1 _102_ (.A(net9),
    .B(_039_),
    .C(_042_),
    .Y(_045_));
 sky130_fd_sc_hd__xnor2_1 _103_ (.A(net10),
    .B(_045_),
    .Y(_005_));
 sky130_fd_sc_hd__xor2_1 _104_ (.A(_068_),
    .B(net12),
    .X(_006_));
 sky130_fd_sc_hd__xor2_1 _105_ (.A(_070_),
    .B(net15),
    .X(_007_));
 sky130_fd_sc_hd__xor2_1 _106_ (.A(_072_),
    .B(net17),
    .X(_008_));
 sky130_fd_sc_hd__nand4_1 _107_ (.A(net9),
    .B(net10),
    .C(net12),
    .D(net11),
    .Y(_020_));
 sky130_fd_sc_hd__nand2_1 _108_ (.A(net15),
    .B(net14),
    .Y(_021_));
 sky130_fd_sc_hd__nor2_1 _109_ (.A(_020_),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__nand3_1 _110_ (.A(net17),
    .B(net16),
    .C(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_1 _111_ (.A(_044_),
    .B(_023_),
    .Y(_073_));
 sky130_fd_sc_hd__xor2_1 _112_ (.A(_074_),
    .B(net19),
    .X(_009_));
 sky130_fd_sc_hd__xor2_1 _113_ (.A(_076_),
    .B(net21),
    .X(_010_));
 sky130_fd_sc_hd__nand2_1 _114_ (.A(net17),
    .B(net16),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _115_ (.A(net19),
    .B(net18),
    .Y(_025_));
 sky130_fd_sc_hd__nand2_1 _116_ (.A(net21),
    .B(net20),
    .Y(_026_));
 sky130_fd_sc_hd__nor3_1 _117_ (.A(_024_),
    .B(_025_),
    .C(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__nand4_1 _118_ (.A(_042_),
    .B(_043_),
    .C(_022_),
    .D(_027_),
    .Y(_028_));
 sky130_fd_sc_hd__xnor2_1 _119_ (.A(net22),
    .B(_028_),
    .Y(_011_));
 sky130_fd_sc_hd__inv_12 _120_ (.A(net1),
    .Y(_019_));
 sky130_fd_sc_hd__nand2_1 _121_ (.A(net25),
    .B(net26),
    .Y(_029_));
 sky130_fd_sc_hd__nor2_1 _122_ (.A(_038_),
    .B(_029_),
    .Y(_059_));
 sky130_fd_sc_hd__and2_0 _123_ (.A(net30),
    .B(_039_),
    .X(_061_));
 sky130_fd_sc_hd__nor4_1 _124_ (.A(_035_),
    .B(_038_),
    .C(_036_),
    .D(_041_),
    .Y(_063_));
 sky130_fd_sc_hd__and3_1 _125_ (.A(net6),
    .B(net5),
    .C(_063_),
    .X(_065_));
 sky130_fd_sc_hd__nand2_1 _126_ (.A(net9),
    .B(net10),
    .Y(_030_));
 sky130_fd_sc_hd__nand2_1 _127_ (.A(_039_),
    .B(_042_),
    .Y(_031_));
 sky130_fd_sc_hd__nor2_1 _128_ (.A(_030_),
    .B(_031_),
    .Y(_067_));
 sky130_fd_sc_hd__nor2_1 _129_ (.A(_020_),
    .B(_031_),
    .Y(_069_));
 sky130_fd_sc_hd__nor3_1 _130_ (.A(_020_),
    .B(_021_),
    .C(_031_),
    .Y(_071_));
 sky130_fd_sc_hd__nor3_1 _131_ (.A(_044_),
    .B(_023_),
    .C(_025_),
    .Y(_075_));
 sky130_fd_sc_hd__ha_1 _132_ (.A(net2),
    .B(net13),
    .COUT(_056_),
    .SUM(_050_));
 sky130_fd_sc_hd__ha_1 _133_ (.A(net2),
    .B(net13),
    .COUT(_057_),
    .SUM(_058_));
 sky130_fd_sc_hd__ha_1 _134_ (.A(net27),
    .B(_059_),
    .COUT(_060_),
    .SUM(_055_));
 sky130_fd_sc_hd__ha_1 _135_ (.A(net3),
    .B(_061_),
    .COUT(_062_),
    .SUM(_046_));
 sky130_fd_sc_hd__ha_1 _136_ (.A(net5),
    .B(_063_),
    .COUT(_064_),
    .SUM(_047_));
 sky130_fd_sc_hd__ha_1 _137_ (.A(net7),
    .B(_065_),
    .COUT(_066_),
    .SUM(_048_));
 sky130_fd_sc_hd__ha_1 _138_ (.A(net11),
    .B(_067_),
    .COUT(_068_),
    .SUM(_049_));
 sky130_fd_sc_hd__ha_1 _139_ (.A(net14),
    .B(_069_),
    .COUT(_070_),
    .SUM(_051_));
 sky130_fd_sc_hd__ha_1 _140_ (.A(net16),
    .B(_071_),
    .COUT(_072_),
    .SUM(_052_));
 sky130_fd_sc_hd__ha_1 _141_ (.A(net18),
    .B(_073_),
    .COUT(_074_),
    .SUM(_053_));
 sky130_fd_sc_hd__ha_1 _142_ (.A(net20),
    .B(_075_),
    .COUT(_076_),
    .SUM(_054_));
 sky130_fd_sc_hd__dfrtp_1 _143_ (.D(_003_),
    .Q(net8),
    .RESET_B(_019_),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.D(_004_),
    .Q(net9),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _145_ (.D(_005_),
    .Q(net10),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _146_ (.D(_049_),
    .Q(net11),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _147_ (.D(_006_),
    .Q(net12),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _148_ (.D(_051_),
    .Q(net14),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _149_ (.D(_007_),
    .Q(net15),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _150_ (.D(_052_),
    .Q(net16),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _151_ (.D(_008_),
    .Q(net17),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _152_ (.D(_053_),
    .Q(net18),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _153_ (.D(_009_),
    .Q(net19),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _154_ (.D(_054_),
    .Q(net20),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _155_ (.D(_010_),
    .Q(net21),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _156_ (.D(_011_),
    .Q(net22),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _157_ (.D(_000_),
    .Q(net2),
    .RESET_B(_019_),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _158_ (.D(_050_),
    .Q(net13),
    .RESET_B(_019_),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 _159_ (.D(_012_),
    .Q(net23),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _160_ (.D(_013_),
    .Q(net24),
    .RESET_B(_019_),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 _161_ (.D(_014_),
    .Q(net25),
    .RESET_B(_019_),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _162_ (.D(_015_),
    .Q(net26),
    .RESET_B(_019_),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _163_ (.D(_055_),
    .Q(net27),
    .RESET_B(_019_),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _164_ (.D(_016_),
    .Q(net28),
    .RESET_B(_019_),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _165_ (.D(_017_),
    .Q(net29),
    .RESET_B(_019_),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _166_ (.D(_018_),
    .Q(net30),
    .RESET_B(_019_),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _167_ (.D(_046_),
    .Q(net3),
    .RESET_B(_019_),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _168_ (.D(_001_),
    .Q(net4),
    .RESET_B(_019_),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _169_ (.D(_047_),
    .Q(net5),
    .RESET_B(_019_),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _170_ (.D(_002_),
    .Q(net6),
    .RESET_B(_019_),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _171_ (.D(_048_),
    .Q(net7),
    .RESET_B(_019_),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_15 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 output2 (.A(net2),
    .X(out[0]));
 sky130_fd_sc_hd__clkbuf_1 output3 (.A(net3),
    .X(out[10]));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net4),
    .X(out[11]));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net5),
    .X(out[12]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net6),
    .X(out[13]));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net7),
    .X(out[14]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net8),
    .X(out[15]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net9),
    .X(out[16]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(out[17]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(out[18]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net12),
    .X(out[19]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .X(out[1]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(out[20]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(out[21]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(out[22]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(out[23]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(out[24]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(out[25]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(out[26]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(out[27]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(out[28]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(out[2]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(out[3]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(out[4]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(out[5]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(out[6]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(out[7]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(out[8]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(out[9]));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_7_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_81 ();
endmodule
